library ieee;
use ieee.std_logic_1164.all;
entity aissa is
 port (
        fom : in std_logic;
        khcham : out std_logic
 );
 end entity;
 